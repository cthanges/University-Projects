----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    15:00:29 10/30/2024 
-- Design Name: 
-- Module Name:    hPosCounter - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity hPosCounter is
    Port ( 
		clk : in  STD_LOGIC);
end hPosCounter;

architecture Behavioral of hPosCounter is

begin
--on clk
--if HD+HFP+HSP+HSB=639
--hpos<= 0
--else: hpos<= hpos+1


end Behavioral;

